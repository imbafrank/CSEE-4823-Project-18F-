

// *********************************************************************************
// Project Name : CSEE 4823 Project: Neural Network Accelerator
// File Name    : nn.v
// Module Name  : nn
// *********************************************************************************
// Modification History:
// Date         By              Version                 Change Description
// -----------------------------------------------------------------------
// 11/13/2018 Shixin Qin      1.0                     Basic function design
// 
// *********************************************************************************

module nn (clk, rst);
    input               clk, rst ;

/*Contol Signal*/
//(for each) memory 

//alu 
	wire alu_op

//agg 


/*Instantiate Module*/


//(for each) memory 

//alu 
	alu ist_alu(
		.rst(rst),  
		(alu_in_a_lsb), 
		(alu_in_b), 
		(alu_op),
		(alu_out)
);

//agg 






endmodule