`include "ctrl_signal.v"

// *********************************************************************************
// Project Name : CSEE 4823 Project: Neural Network Accelerator
// File Name    : ctrl.v
// *********************************************************************************
// Modification History:
// Date         By              Version                 Change Description
// -----------------------------------------------------------------------
// 11/13/2018 	Shixin Qin      1.0                     Basic function design
// 
// *********************************************************************************

module ctrl (clk, rst,  );
    input               clk, rst ;
    output               ;

    always @()
    begin

    end
endmodule